module xml

pub const header = '<?xml version="1.0" encoding="utf-8"?>'
